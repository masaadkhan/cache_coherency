module top ();

  cache c1 ();
  cache c2 ();
  cache c3 ();

endmodule
